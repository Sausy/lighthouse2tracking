
module PolyFinder (
      input  [16:0] io_startState,
      input  [16:0] io_targetState,
      input  [9:0] io_maxTick,
      input   io_start_valid,
      output  io_start_ready,
      output  io_found,
      output [4:0] io_polyFound,
      output  io_done_valid,
      input   io_done_ready,
      input   Slow_clk);
  wire  _zz_96_;
  wire  _zz_97_;
  wire  _zz_98_;
  wire  _zz_99_;
  wire  _zz_100_;
  wire  _zz_101_;
  wire  _zz_102_;
  wire  _zz_103_;
  wire  _zz_104_;
  wire  _zz_105_;
  wire  _zz_106_;
  wire  _zz_107_;
  wire  _zz_108_;
  wire  _zz_109_;
  wire  _zz_110_;
  wire  _zz_111_;
  wire  _zz_112_;
  wire  _zz_113_;
  wire  _zz_114_;
  wire  _zz_115_;
  wire  _zz_116_;
  wire  _zz_117_;
  wire  _zz_118_;
  wire  _zz_119_;
  wire  _zz_120_;
  wire  _zz_121_;
  wire  _zz_122_;
  wire  _zz_123_;
  wire  _zz_124_;
  wire  _zz_125_;
  wire  _zz_126_;
  wire  _zz_127_;
  wire  _zz_128_;
  wire  _zz_129_;
  wire  _zz_130_;
  wire  _zz_131_;
  wire  _zz_132_;
  wire  _zz_133_;
  wire  _zz_134_;
  wire  _zz_135_;
  wire  _zz_136_;
  wire  _zz_137_;
  wire  _zz_138_;
  wire  _zz_139_;
  wire  _zz_140_;
  wire  _zz_141_;
  wire  _zz_142_;
  wire  _zz_143_;
  wire  _zz_144_;
  wire  _zz_145_;
  wire  _zz_146_;
  wire  _zz_147_;
  wire  _zz_148_;
  wire  _zz_149_;
  wire  _zz_150_;
  wire  _zz_151_;
  wire  _zz_152_;
  wire  _zz_153_;
  wire  _zz_154_;
  wire  _zz_155_;
  wire  _zz_156_;
  wire  _zz_157_;
  wire  _zz_158_;
  wire  _zz_159_;
  reg  searching = 1'b0;
  reg [31:0] found = (32'b00000000000000000000000000000000);
  wire  _zz_1_;
  wire  _zz_2_;
  wire  _zz_3_;
  wire  _zz_4_;
  wire  _zz_5_;
  wire  _zz_6_;
  wire  _zz_7_;
  wire  _zz_8_;
  wire  _zz_9_;
  wire  _zz_10_;
  wire  _zz_11_;
  wire  _zz_12_;
  wire  _zz_13_;
  wire  _zz_14_;
  wire  _zz_15_;
  wire  _zz_16_;
  wire  _zz_17_;
  wire  _zz_18_;
  wire  _zz_19_;
  wire  _zz_20_;
  wire  _zz_21_;
  wire  _zz_22_;
  wire  _zz_23_;
  wire  _zz_24_;
  wire  _zz_25_;
  wire  _zz_26_;
  wire  _zz_27_;
  wire  _zz_28_;
  wire  _zz_29_;
  wire  _zz_30_;
  wire  _zz_31_;
  reg  searching_regNext;
  reg [9:0] counter = (10'b0000000000);
  wire [16:0] states_0;
  wire [16:0] states_1;
  wire [16:0] states_2;
  wire [16:0] states_3;
  wire [16:0] states_4;
  wire [16:0] states_5;
  wire [16:0] states_6;
  wire [16:0] states_7;
  wire [16:0] states_8;
  wire [16:0] states_9;
  wire [16:0] states_10;
  wire [16:0] states_11;
  wire [16:0] states_12;
  wire [16:0] states_13;
  wire [16:0] states_14;
  wire [16:0] states_15;
  wire [16:0] states_16;
  wire [16:0] states_17;
  wire [16:0] states_18;
  wire [16:0] states_19;
  wire [16:0] states_20;
  wire [16:0] states_21;
  wire [16:0] states_22;
  wire [16:0] states_23;
  wire [16:0] states_24;
  wire [16:0] states_25;
  wire [16:0] states_26;
  wire [16:0] states_27;
  wire [16:0] states_28;
  wire [16:0] states_29;
  wire [16:0] states_30;
  wire [16:0] states_31;
  reg [16:0] _zz_32_ = (17'b00000000000000000);
  wire [16:0] _zz_33_;
  reg [16:0] _zz_34_ = (17'b00000000000000000);
  wire [16:0] _zz_35_;
  reg [16:0] _zz_36_ = (17'b00000000000000000);
  wire [16:0] _zz_37_;
  reg [16:0] _zz_38_ = (17'b00000000000000000);
  wire [16:0] _zz_39_;
  reg [16:0] _zz_40_ = (17'b00000000000000000);
  wire [16:0] _zz_41_;
  reg [16:0] _zz_42_ = (17'b00000000000000000);
  wire [16:0] _zz_43_;
  reg [16:0] _zz_44_ = (17'b00000000000000000);
  wire [16:0] _zz_45_;
  reg [16:0] _zz_46_ = (17'b00000000000000000);
  wire [16:0] _zz_47_;
  reg [16:0] _zz_48_ = (17'b00000000000000000);
  wire [16:0] _zz_49_;
  reg [16:0] _zz_50_ = (17'b00000000000000000);
  wire [16:0] _zz_51_;
  reg [16:0] _zz_52_ = (17'b00000000000000000);
  wire [16:0] _zz_53_;
  reg [16:0] _zz_54_ = (17'b00000000000000000);
  wire [16:0] _zz_55_;
  reg [16:0] _zz_56_ = (17'b00000000000000000);
  wire [16:0] _zz_57_;
  reg [16:0] _zz_58_ = (17'b00000000000000000);
  wire [16:0] _zz_59_;
  reg [16:0] _zz_60_ = (17'b00000000000000000);
  wire [16:0] _zz_61_;
  reg [16:0] _zz_62_ = (17'b00000000000000000);
  wire [16:0] _zz_63_;
  reg [16:0] _zz_64_ = (17'b00000000000000000);
  wire [16:0] _zz_65_;
  reg [16:0] _zz_66_ = (17'b00000000000000000);
  wire [16:0] _zz_67_;
  reg [16:0] _zz_68_ = (17'b00000000000000000);
  wire [16:0] _zz_69_;
  reg [16:0] _zz_70_ = (17'b00000000000000000);
  wire [16:0] _zz_71_;
  reg [16:0] _zz_72_ = (17'b00000000000000000);
  wire [16:0] _zz_73_;
  reg [16:0] _zz_74_ = (17'b00000000000000000);
  wire [16:0] _zz_75_;
  reg [16:0] _zz_76_ = (17'b00000000000000000);
  wire [16:0] _zz_77_;
  reg [16:0] _zz_78_ = (17'b00000000000000000);
  wire [16:0] _zz_79_;
  reg [16:0] _zz_80_ = (17'b00000000000000000);
  wire [16:0] _zz_81_;
  reg [16:0] _zz_82_ = (17'b00000000000000000);
  wire [16:0] _zz_83_;
  reg [16:0] _zz_84_ = (17'b00000000000000000);
  wire [16:0] _zz_85_;
  reg [16:0] _zz_86_ = (17'b00000000000000000);
  wire [16:0] _zz_87_;
  reg [16:0] _zz_88_ = (17'b00000000000000000);
  wire [16:0] _zz_89_;
  reg [16:0] _zz_90_ = (17'b00000000000000000);
  wire [16:0] _zz_91_;
  reg [16:0] _zz_92_ = (17'b00000000000000000);
  wire [16:0] _zz_93_;
  reg [16:0] _zz_94_ = (17'b00000000000000000);
  wire [16:0] _zz_95_;
  assign _zz_96_ = ((_zz_33_[0] ^ _zz_33_[1]) ^ _zz_33_[2]);
  assign _zz_97_ = _zz_33_[3];
  assign _zz_98_ = ((_zz_35_[0] ^ _zz_35_[1]) ^ _zz_35_[2]);
  assign _zz_99_ = _zz_35_[3];
  assign _zz_100_ = ((_zz_37_[0] ^ _zz_37_[1]) ^ _zz_37_[2]);
  assign _zz_101_ = _zz_37_[3];
  assign _zz_102_ = ((_zz_39_[0] ^ _zz_39_[1]) ^ _zz_39_[2]);
  assign _zz_103_ = _zz_39_[3];
  assign _zz_104_ = ((_zz_41_[0] ^ _zz_41_[1]) ^ _zz_41_[2]);
  assign _zz_105_ = _zz_41_[3];
  assign _zz_106_ = ((_zz_43_[0] ^ _zz_43_[1]) ^ _zz_43_[2]);
  assign _zz_107_ = _zz_43_[3];
  assign _zz_108_ = ((_zz_45_[0] ^ _zz_45_[1]) ^ _zz_45_[2]);
  assign _zz_109_ = _zz_45_[3];
  assign _zz_110_ = ((_zz_47_[0] ^ _zz_47_[1]) ^ _zz_47_[2]);
  assign _zz_111_ = _zz_47_[3];
  assign _zz_112_ = ((_zz_49_[0] ^ _zz_49_[1]) ^ _zz_49_[2]);
  assign _zz_113_ = _zz_49_[3];
  assign _zz_114_ = ((_zz_51_[0] ^ _zz_51_[1]) ^ _zz_51_[2]);
  assign _zz_115_ = _zz_51_[3];
  assign _zz_116_ = ((_zz_53_[0] ^ _zz_53_[1]) ^ _zz_53_[2]);
  assign _zz_117_ = _zz_53_[3];
  assign _zz_118_ = ((_zz_55_[0] ^ _zz_55_[1]) ^ _zz_55_[2]);
  assign _zz_119_ = _zz_55_[3];
  assign _zz_120_ = ((_zz_57_[0] ^ _zz_57_[1]) ^ _zz_57_[2]);
  assign _zz_121_ = _zz_57_[3];
  assign _zz_122_ = ((_zz_59_[0] ^ _zz_59_[1]) ^ _zz_59_[2]);
  assign _zz_123_ = _zz_59_[3];
  assign _zz_124_ = ((_zz_61_[0] ^ _zz_61_[1]) ^ _zz_61_[2]);
  assign _zz_125_ = _zz_61_[3];
  assign _zz_126_ = ((_zz_63_[0] ^ _zz_63_[1]) ^ _zz_63_[2]);
  assign _zz_127_ = _zz_63_[3];
  assign _zz_128_ = ((_zz_65_[0] ^ _zz_65_[1]) ^ _zz_65_[2]);
  assign _zz_129_ = _zz_65_[3];
  assign _zz_130_ = ((_zz_67_[0] ^ _zz_67_[1]) ^ _zz_67_[2]);
  assign _zz_131_ = _zz_67_[3];
  assign _zz_132_ = ((_zz_69_[0] ^ _zz_69_[1]) ^ _zz_69_[2]);
  assign _zz_133_ = _zz_69_[3];
  assign _zz_134_ = ((_zz_71_[0] ^ _zz_71_[1]) ^ _zz_71_[2]);
  assign _zz_135_ = _zz_71_[3];
  assign _zz_136_ = ((_zz_73_[0] ^ _zz_73_[1]) ^ _zz_73_[2]);
  assign _zz_137_ = _zz_73_[3];
  assign _zz_138_ = ((_zz_75_[0] ^ _zz_75_[1]) ^ _zz_75_[2]);
  assign _zz_139_ = _zz_75_[3];
  assign _zz_140_ = ((_zz_77_[0] ^ _zz_77_[1]) ^ _zz_77_[2]);
  assign _zz_141_ = _zz_77_[3];
  assign _zz_142_ = ((_zz_79_[0] ^ _zz_79_[1]) ^ _zz_79_[2]);
  assign _zz_143_ = _zz_79_[3];
  assign _zz_144_ = ((_zz_81_[0] ^ _zz_81_[1]) ^ _zz_81_[2]);
  assign _zz_145_ = _zz_81_[3];
  assign _zz_146_ = ((_zz_83_[0] ^ _zz_83_[1]) ^ _zz_83_[2]);
  assign _zz_147_ = _zz_83_[3];
  assign _zz_148_ = ((_zz_85_[0] ^ _zz_85_[1]) ^ _zz_85_[2]);
  assign _zz_149_ = _zz_85_[3];
  assign _zz_150_ = ((_zz_87_[0] ^ _zz_87_[1]) ^ _zz_87_[2]);
  assign _zz_151_ = _zz_87_[3];
  assign _zz_152_ = ((_zz_89_[0] ^ _zz_89_[1]) ^ _zz_89_[2]);
  assign _zz_153_ = _zz_89_[3];
  assign _zz_154_ = ((_zz_91_[0] ^ _zz_91_[1]) ^ _zz_91_[2]);
  assign _zz_155_ = _zz_91_[3];
  assign _zz_156_ = ((_zz_93_[0] ^ _zz_93_[1]) ^ _zz_93_[2]);
  assign _zz_157_ = _zz_93_[3];
  assign _zz_158_ = ((_zz_95_[0] ^ _zz_95_[1]) ^ _zz_95_[2]);
  assign _zz_159_ = _zz_95_[3];
  assign _zz_1_ = found[3];
  assign _zz_2_ = found[5];
  assign _zz_3_ = found[6];
  assign _zz_4_ = found[7];
  assign _zz_5_ = found[9];
  assign _zz_6_ = found[10];
  assign _zz_7_ = found[11];
  assign _zz_8_ = found[12];
  assign _zz_9_ = found[13];
  assign _zz_10_ = found[14];
  assign _zz_11_ = found[15];
  assign _zz_12_ = found[17];
  assign _zz_13_ = found[18];
  assign _zz_14_ = found[19];
  assign _zz_15_ = found[20];
  assign _zz_16_ = found[21];
  assign _zz_17_ = found[22];
  assign _zz_18_ = found[23];
  assign _zz_19_ = found[24];
  assign _zz_20_ = found[25];
  assign _zz_21_ = found[26];
  assign _zz_22_ = found[27];
  assign _zz_23_ = found[28];
  assign _zz_24_ = found[29];
  assign _zz_25_ = found[30];
  assign _zz_26_ = found[31];
  assign _zz_27_ = (((((((((((((((found[1] || _zz_1_) || _zz_2_) || _zz_4_) || _zz_5_) || _zz_7_) || _zz_9_) || _zz_11_) || _zz_12_) || _zz_14_) || _zz_16_) || _zz_18_) || _zz_20_) || _zz_22_) || _zz_24_) || _zz_26_);
  assign _zz_28_ = (((((((((((((((found[2] || _zz_1_) || _zz_3_) || _zz_4_) || _zz_6_) || _zz_7_) || _zz_10_) || _zz_11_) || _zz_13_) || _zz_14_) || _zz_17_) || _zz_18_) || _zz_21_) || _zz_22_) || _zz_25_) || _zz_26_);
  assign _zz_29_ = (((((((((((((((found[4] || _zz_2_) || _zz_3_) || _zz_4_) || _zz_8_) || _zz_9_) || _zz_10_) || _zz_11_) || _zz_15_) || _zz_16_) || _zz_17_) || _zz_18_) || _zz_23_) || _zz_24_) || _zz_25_) || _zz_26_);
  assign _zz_30_ = (((((((((((((((found[8] || _zz_5_) || _zz_6_) || _zz_7_) || _zz_8_) || _zz_9_) || _zz_10_) || _zz_11_) || _zz_19_) || _zz_20_) || _zz_21_) || _zz_22_) || _zz_23_) || _zz_24_) || _zz_25_) || _zz_26_);
  assign _zz_31_ = (((((((((((((((found[16] || _zz_12_) || _zz_13_) || _zz_14_) || _zz_15_) || _zz_16_) || _zz_17_) || _zz_18_) || _zz_19_) || _zz_20_) || _zz_21_) || _zz_22_) || _zz_23_) || _zz_24_) || _zz_25_) || _zz_26_);
  assign io_polyFound = {_zz_31_,{_zz_30_,{_zz_29_,{_zz_28_,_zz_27_}}}};
  assign io_done_valid = ((! searching) && searching_regNext);
  assign io_found = (found != (32'b00000000000000000000000000000000));
  assign io_start_ready = 1'b1;
  assign states_0 = _zz_32_;
  assign _zz_33_ = (_zz_32_ & (17'b11101001001011000));
  assign states_1 = _zz_34_;
  assign _zz_35_ = (_zz_34_ & (17'b10111111000000100));
  assign states_2 = _zz_36_;
  assign _zz_37_ = (_zz_36_ & (17'b11111111101101011));
  assign states_3 = _zz_38_;
  assign _zz_39_ = (_zz_38_ & (17'b10011111101100111));
  assign states_4 = _zz_40_;
  assign _zz_41_ = (_zz_40_ & (17'b11011100111101110));
  assign states_5 = _zz_42_;
  assign _zz_43_ = (_zz_42_ & (17'b11001100011010001));
  assign states_6 = _zz_44_;
  assign _zz_45_ = (_zz_44_ & (17'b10111100011000111));
  assign states_7 = _zz_46_;
  assign _zz_47_ = (_zz_46_ & (17'b11000101001010101));
  assign states_8 = _zz_48_;
  assign _zz_49_ = (_zz_48_ & (17'b10101011101110111));
  assign states_9 = _zz_50_;
  assign _zz_51_ = (_zz_50_ & (17'b11101100100010001));
  assign states_10 = _zz_52_;
  assign _zz_53_ = (_zz_52_ & (17'b10101011101101001));
  assign states_11 = _zz_54_;
  assign _zz_55_ = (_zz_54_ & (17'b11001100100011111));
  assign states_12 = _zz_56_;
  assign _zz_57_ = (_zz_56_ & (17'b10010101111010000));
  assign states_13 = _zz_58_;
  assign _zz_59_ = (_zz_58_ & (17'b11100111101110011));
  assign states_14 = _zz_60_;
  assign _zz_61_ = (_zz_60_ & (17'b10011011001011101));
  assign states_15 = _zz_62_;
  assign _zz_63_ = (_zz_62_ & (17'b11001011111110101));
  assign states_16 = _zz_64_;
  assign _zz_65_ = (_zz_64_ & (17'b11001010010100000));
  assign states_17 = _zz_66_;
  assign _zz_67_ = (_zz_66_ & (17'b11011001001111001));
  assign states_18 = _zz_68_;
  assign _zz_69_ = (_zz_68_ & (17'b10011101000110100));
  assign states_19 = _zz_70_;
  assign _zz_71_ = (_zz_70_ & (17'b11010111001000001));
  assign states_20 = _zz_72_;
  assign _zz_73_ = (_zz_72_ & (17'b11000000011010100));
  assign states_21 = _zz_74_;
  assign _zz_75_ = (_zz_74_ & (17'b10111100010010001));
  assign states_22 = _zz_76_;
  assign _zz_77_ = (_zz_76_ & (17'b10010111001100100));
  assign states_23 = _zz_78_;
  assign _zz_79_ = (_zz_78_ & (17'b10111110001110010));
  assign states_24 = _zz_80_;
  assign _zz_81_ = (_zz_80_ & (17'b11001110001101101));
  assign states_25 = _zz_82_;
  assign _zz_83_ = (_zz_82_ & (17'b10011111100110010));
  assign states_26 = _zz_84_;
  assign _zz_85_ = (_zz_84_ & (17'b11010111000010100));
  assign states_27 = _zz_86_;
  assign _zz_87_ = (_zz_86_ & (17'b10100111001110110));
  assign states_28 = _zz_88_;
  assign _zz_89_ = (_zz_88_ & (17'b10011110010010111));
  assign states_29 = _zz_90_;
  assign _zz_91_ = (_zz_90_ & (17'b10011000011001011));
  assign states_30 = _zz_92_;
  assign _zz_93_ = (_zz_92_ & (17'b10011011101010000));
  assign states_31 = _zz_94_;
  assign _zz_95_ = (_zz_94_ & (17'b11100101110001101));
  always @ (posedge Slow_clk) begin
    if(searching)begin
      counter <= (counter - (10'b0000000001));
      if((counter == (10'b0000000000)))begin
        searching <= 1'b0;
        found <= (32'b00000000000000000000000000000000);
      end
    end else begin
      counter <= io_maxTick;
    end
    if((io_start_valid && io_start_ready))begin
      searching <= 1'b1;
      found <= (32'b00000000000000000000000000000000);
    end
    if((io_start_valid && io_start_ready))begin
      _zz_32_ <= io_startState;
    end
    if(searching)begin
      _zz_32_ <= {_zz_32_[15 : 0],((((((((((((((_zz_96_ ^ _zz_97_) ^ _zz_33_[4]) ^ _zz_33_[5]) ^ _zz_33_[6]) ^ _zz_33_[7]) ^ _zz_33_[8]) ^ _zz_33_[9]) ^ _zz_33_[10]) ^ _zz_33_[11]) ^ _zz_33_[12]) ^ _zz_33_[13]) ^ _zz_33_[14]) ^ _zz_33_[15]) ^ _zz_33_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_32_ == io_targetState)))begin
        found[0] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_34_ <= io_startState;
    end
    if(searching)begin
      _zz_34_ <= {_zz_34_[15 : 0],((((((((((((((_zz_98_ ^ _zz_99_) ^ _zz_35_[4]) ^ _zz_35_[5]) ^ _zz_35_[6]) ^ _zz_35_[7]) ^ _zz_35_[8]) ^ _zz_35_[9]) ^ _zz_35_[10]) ^ _zz_35_[11]) ^ _zz_35_[12]) ^ _zz_35_[13]) ^ _zz_35_[14]) ^ _zz_35_[15]) ^ _zz_35_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_34_ == io_targetState)))begin
        found[1] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_36_ <= io_startState;
    end
    if(searching)begin
      _zz_36_ <= {_zz_36_[15 : 0],((((((((((((((_zz_100_ ^ _zz_101_) ^ _zz_37_[4]) ^ _zz_37_[5]) ^ _zz_37_[6]) ^ _zz_37_[7]) ^ _zz_37_[8]) ^ _zz_37_[9]) ^ _zz_37_[10]) ^ _zz_37_[11]) ^ _zz_37_[12]) ^ _zz_37_[13]) ^ _zz_37_[14]) ^ _zz_37_[15]) ^ _zz_37_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_36_ == io_targetState)))begin
        found[2] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_38_ <= io_startState;
    end
    if(searching)begin
      _zz_38_ <= {_zz_38_[15 : 0],((((((((((((((_zz_102_ ^ _zz_103_) ^ _zz_39_[4]) ^ _zz_39_[5]) ^ _zz_39_[6]) ^ _zz_39_[7]) ^ _zz_39_[8]) ^ _zz_39_[9]) ^ _zz_39_[10]) ^ _zz_39_[11]) ^ _zz_39_[12]) ^ _zz_39_[13]) ^ _zz_39_[14]) ^ _zz_39_[15]) ^ _zz_39_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_38_ == io_targetState)))begin
        found[3] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_40_ <= io_startState;
    end
    if(searching)begin
      _zz_40_ <= {_zz_40_[15 : 0],((((((((((((((_zz_104_ ^ _zz_105_) ^ _zz_41_[4]) ^ _zz_41_[5]) ^ _zz_41_[6]) ^ _zz_41_[7]) ^ _zz_41_[8]) ^ _zz_41_[9]) ^ _zz_41_[10]) ^ _zz_41_[11]) ^ _zz_41_[12]) ^ _zz_41_[13]) ^ _zz_41_[14]) ^ _zz_41_[15]) ^ _zz_41_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_40_ == io_targetState)))begin
        found[4] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_42_ <= io_startState;
    end
    if(searching)begin
      _zz_42_ <= {_zz_42_[15 : 0],((((((((((((((_zz_106_ ^ _zz_107_) ^ _zz_43_[4]) ^ _zz_43_[5]) ^ _zz_43_[6]) ^ _zz_43_[7]) ^ _zz_43_[8]) ^ _zz_43_[9]) ^ _zz_43_[10]) ^ _zz_43_[11]) ^ _zz_43_[12]) ^ _zz_43_[13]) ^ _zz_43_[14]) ^ _zz_43_[15]) ^ _zz_43_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_42_ == io_targetState)))begin
        found[5] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_44_ <= io_startState;
    end
    if(searching)begin
      _zz_44_ <= {_zz_44_[15 : 0],((((((((((((((_zz_108_ ^ _zz_109_) ^ _zz_45_[4]) ^ _zz_45_[5]) ^ _zz_45_[6]) ^ _zz_45_[7]) ^ _zz_45_[8]) ^ _zz_45_[9]) ^ _zz_45_[10]) ^ _zz_45_[11]) ^ _zz_45_[12]) ^ _zz_45_[13]) ^ _zz_45_[14]) ^ _zz_45_[15]) ^ _zz_45_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_44_ == io_targetState)))begin
        found[6] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_46_ <= io_startState;
    end
    if(searching)begin
      _zz_46_ <= {_zz_46_[15 : 0],((((((((((((((_zz_110_ ^ _zz_111_) ^ _zz_47_[4]) ^ _zz_47_[5]) ^ _zz_47_[6]) ^ _zz_47_[7]) ^ _zz_47_[8]) ^ _zz_47_[9]) ^ _zz_47_[10]) ^ _zz_47_[11]) ^ _zz_47_[12]) ^ _zz_47_[13]) ^ _zz_47_[14]) ^ _zz_47_[15]) ^ _zz_47_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_46_ == io_targetState)))begin
        found[7] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_48_ <= io_startState;
    end
    if(searching)begin
      _zz_48_ <= {_zz_48_[15 : 0],((((((((((((((_zz_112_ ^ _zz_113_) ^ _zz_49_[4]) ^ _zz_49_[5]) ^ _zz_49_[6]) ^ _zz_49_[7]) ^ _zz_49_[8]) ^ _zz_49_[9]) ^ _zz_49_[10]) ^ _zz_49_[11]) ^ _zz_49_[12]) ^ _zz_49_[13]) ^ _zz_49_[14]) ^ _zz_49_[15]) ^ _zz_49_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_48_ == io_targetState)))begin
        found[8] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_50_ <= io_startState;
    end
    if(searching)begin
      _zz_50_ <= {_zz_50_[15 : 0],((((((((((((((_zz_114_ ^ _zz_115_) ^ _zz_51_[4]) ^ _zz_51_[5]) ^ _zz_51_[6]) ^ _zz_51_[7]) ^ _zz_51_[8]) ^ _zz_51_[9]) ^ _zz_51_[10]) ^ _zz_51_[11]) ^ _zz_51_[12]) ^ _zz_51_[13]) ^ _zz_51_[14]) ^ _zz_51_[15]) ^ _zz_51_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_50_ == io_targetState)))begin
        found[9] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_52_ <= io_startState;
    end
    if(searching)begin
      _zz_52_ <= {_zz_52_[15 : 0],((((((((((((((_zz_116_ ^ _zz_117_) ^ _zz_53_[4]) ^ _zz_53_[5]) ^ _zz_53_[6]) ^ _zz_53_[7]) ^ _zz_53_[8]) ^ _zz_53_[9]) ^ _zz_53_[10]) ^ _zz_53_[11]) ^ _zz_53_[12]) ^ _zz_53_[13]) ^ _zz_53_[14]) ^ _zz_53_[15]) ^ _zz_53_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_52_ == io_targetState)))begin
        found[10] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_54_ <= io_startState;
    end
    if(searching)begin
      _zz_54_ <= {_zz_54_[15 : 0],((((((((((((((_zz_118_ ^ _zz_119_) ^ _zz_55_[4]) ^ _zz_55_[5]) ^ _zz_55_[6]) ^ _zz_55_[7]) ^ _zz_55_[8]) ^ _zz_55_[9]) ^ _zz_55_[10]) ^ _zz_55_[11]) ^ _zz_55_[12]) ^ _zz_55_[13]) ^ _zz_55_[14]) ^ _zz_55_[15]) ^ _zz_55_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_54_ == io_targetState)))begin
        found[11] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_56_ <= io_startState;
    end
    if(searching)begin
      _zz_56_ <= {_zz_56_[15 : 0],((((((((((((((_zz_120_ ^ _zz_121_) ^ _zz_57_[4]) ^ _zz_57_[5]) ^ _zz_57_[6]) ^ _zz_57_[7]) ^ _zz_57_[8]) ^ _zz_57_[9]) ^ _zz_57_[10]) ^ _zz_57_[11]) ^ _zz_57_[12]) ^ _zz_57_[13]) ^ _zz_57_[14]) ^ _zz_57_[15]) ^ _zz_57_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_56_ == io_targetState)))begin
        found[12] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_58_ <= io_startState;
    end
    if(searching)begin
      _zz_58_ <= {_zz_58_[15 : 0],((((((((((((((_zz_122_ ^ _zz_123_) ^ _zz_59_[4]) ^ _zz_59_[5]) ^ _zz_59_[6]) ^ _zz_59_[7]) ^ _zz_59_[8]) ^ _zz_59_[9]) ^ _zz_59_[10]) ^ _zz_59_[11]) ^ _zz_59_[12]) ^ _zz_59_[13]) ^ _zz_59_[14]) ^ _zz_59_[15]) ^ _zz_59_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_58_ == io_targetState)))begin
        found[13] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_60_ <= io_startState;
    end
    if(searching)begin
      _zz_60_ <= {_zz_60_[15 : 0],((((((((((((((_zz_124_ ^ _zz_125_) ^ _zz_61_[4]) ^ _zz_61_[5]) ^ _zz_61_[6]) ^ _zz_61_[7]) ^ _zz_61_[8]) ^ _zz_61_[9]) ^ _zz_61_[10]) ^ _zz_61_[11]) ^ _zz_61_[12]) ^ _zz_61_[13]) ^ _zz_61_[14]) ^ _zz_61_[15]) ^ _zz_61_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_60_ == io_targetState)))begin
        found[14] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_62_ <= io_startState;
    end
    if(searching)begin
      _zz_62_ <= {_zz_62_[15 : 0],((((((((((((((_zz_126_ ^ _zz_127_) ^ _zz_63_[4]) ^ _zz_63_[5]) ^ _zz_63_[6]) ^ _zz_63_[7]) ^ _zz_63_[8]) ^ _zz_63_[9]) ^ _zz_63_[10]) ^ _zz_63_[11]) ^ _zz_63_[12]) ^ _zz_63_[13]) ^ _zz_63_[14]) ^ _zz_63_[15]) ^ _zz_63_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_62_ == io_targetState)))begin
        found[15] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_64_ <= io_startState;
    end
    if(searching)begin
      _zz_64_ <= {_zz_64_[15 : 0],((((((((((((((_zz_128_ ^ _zz_129_) ^ _zz_65_[4]) ^ _zz_65_[5]) ^ _zz_65_[6]) ^ _zz_65_[7]) ^ _zz_65_[8]) ^ _zz_65_[9]) ^ _zz_65_[10]) ^ _zz_65_[11]) ^ _zz_65_[12]) ^ _zz_65_[13]) ^ _zz_65_[14]) ^ _zz_65_[15]) ^ _zz_65_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_64_ == io_targetState)))begin
        found[16] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_66_ <= io_startState;
    end
    if(searching)begin
      _zz_66_ <= {_zz_66_[15 : 0],((((((((((((((_zz_130_ ^ _zz_131_) ^ _zz_67_[4]) ^ _zz_67_[5]) ^ _zz_67_[6]) ^ _zz_67_[7]) ^ _zz_67_[8]) ^ _zz_67_[9]) ^ _zz_67_[10]) ^ _zz_67_[11]) ^ _zz_67_[12]) ^ _zz_67_[13]) ^ _zz_67_[14]) ^ _zz_67_[15]) ^ _zz_67_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_66_ == io_targetState)))begin
        found[17] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_68_ <= io_startState;
    end
    if(searching)begin
      _zz_68_ <= {_zz_68_[15 : 0],((((((((((((((_zz_132_ ^ _zz_133_) ^ _zz_69_[4]) ^ _zz_69_[5]) ^ _zz_69_[6]) ^ _zz_69_[7]) ^ _zz_69_[8]) ^ _zz_69_[9]) ^ _zz_69_[10]) ^ _zz_69_[11]) ^ _zz_69_[12]) ^ _zz_69_[13]) ^ _zz_69_[14]) ^ _zz_69_[15]) ^ _zz_69_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_68_ == io_targetState)))begin
        found[18] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_70_ <= io_startState;
    end
    if(searching)begin
      _zz_70_ <= {_zz_70_[15 : 0],((((((((((((((_zz_134_ ^ _zz_135_) ^ _zz_71_[4]) ^ _zz_71_[5]) ^ _zz_71_[6]) ^ _zz_71_[7]) ^ _zz_71_[8]) ^ _zz_71_[9]) ^ _zz_71_[10]) ^ _zz_71_[11]) ^ _zz_71_[12]) ^ _zz_71_[13]) ^ _zz_71_[14]) ^ _zz_71_[15]) ^ _zz_71_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_70_ == io_targetState)))begin
        found[19] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_72_ <= io_startState;
    end
    if(searching)begin
      _zz_72_ <= {_zz_72_[15 : 0],((((((((((((((_zz_136_ ^ _zz_137_) ^ _zz_73_[4]) ^ _zz_73_[5]) ^ _zz_73_[6]) ^ _zz_73_[7]) ^ _zz_73_[8]) ^ _zz_73_[9]) ^ _zz_73_[10]) ^ _zz_73_[11]) ^ _zz_73_[12]) ^ _zz_73_[13]) ^ _zz_73_[14]) ^ _zz_73_[15]) ^ _zz_73_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_72_ == io_targetState)))begin
        found[20] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_74_ <= io_startState;
    end
    if(searching)begin
      _zz_74_ <= {_zz_74_[15 : 0],((((((((((((((_zz_138_ ^ _zz_139_) ^ _zz_75_[4]) ^ _zz_75_[5]) ^ _zz_75_[6]) ^ _zz_75_[7]) ^ _zz_75_[8]) ^ _zz_75_[9]) ^ _zz_75_[10]) ^ _zz_75_[11]) ^ _zz_75_[12]) ^ _zz_75_[13]) ^ _zz_75_[14]) ^ _zz_75_[15]) ^ _zz_75_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_74_ == io_targetState)))begin
        found[21] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_76_ <= io_startState;
    end
    if(searching)begin
      _zz_76_ <= {_zz_76_[15 : 0],((((((((((((((_zz_140_ ^ _zz_141_) ^ _zz_77_[4]) ^ _zz_77_[5]) ^ _zz_77_[6]) ^ _zz_77_[7]) ^ _zz_77_[8]) ^ _zz_77_[9]) ^ _zz_77_[10]) ^ _zz_77_[11]) ^ _zz_77_[12]) ^ _zz_77_[13]) ^ _zz_77_[14]) ^ _zz_77_[15]) ^ _zz_77_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_76_ == io_targetState)))begin
        found[22] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_78_ <= io_startState;
    end
    if(searching)begin
      _zz_78_ <= {_zz_78_[15 : 0],((((((((((((((_zz_142_ ^ _zz_143_) ^ _zz_79_[4]) ^ _zz_79_[5]) ^ _zz_79_[6]) ^ _zz_79_[7]) ^ _zz_79_[8]) ^ _zz_79_[9]) ^ _zz_79_[10]) ^ _zz_79_[11]) ^ _zz_79_[12]) ^ _zz_79_[13]) ^ _zz_79_[14]) ^ _zz_79_[15]) ^ _zz_79_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_78_ == io_targetState)))begin
        found[23] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_80_ <= io_startState;
    end
    if(searching)begin
      _zz_80_ <= {_zz_80_[15 : 0],((((((((((((((_zz_144_ ^ _zz_145_) ^ _zz_81_[4]) ^ _zz_81_[5]) ^ _zz_81_[6]) ^ _zz_81_[7]) ^ _zz_81_[8]) ^ _zz_81_[9]) ^ _zz_81_[10]) ^ _zz_81_[11]) ^ _zz_81_[12]) ^ _zz_81_[13]) ^ _zz_81_[14]) ^ _zz_81_[15]) ^ _zz_81_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_80_ == io_targetState)))begin
        found[24] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_82_ <= io_startState;
    end
    if(searching)begin
      _zz_82_ <= {_zz_82_[15 : 0],((((((((((((((_zz_146_ ^ _zz_147_) ^ _zz_83_[4]) ^ _zz_83_[5]) ^ _zz_83_[6]) ^ _zz_83_[7]) ^ _zz_83_[8]) ^ _zz_83_[9]) ^ _zz_83_[10]) ^ _zz_83_[11]) ^ _zz_83_[12]) ^ _zz_83_[13]) ^ _zz_83_[14]) ^ _zz_83_[15]) ^ _zz_83_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_82_ == io_targetState)))begin
        found[25] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_84_ <= io_startState;
    end
    if(searching)begin
      _zz_84_ <= {_zz_84_[15 : 0],((((((((((((((_zz_148_ ^ _zz_149_) ^ _zz_85_[4]) ^ _zz_85_[5]) ^ _zz_85_[6]) ^ _zz_85_[7]) ^ _zz_85_[8]) ^ _zz_85_[9]) ^ _zz_85_[10]) ^ _zz_85_[11]) ^ _zz_85_[12]) ^ _zz_85_[13]) ^ _zz_85_[14]) ^ _zz_85_[15]) ^ _zz_85_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_84_ == io_targetState)))begin
        found[26] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_86_ <= io_startState;
    end
    if(searching)begin
      _zz_86_ <= {_zz_86_[15 : 0],((((((((((((((_zz_150_ ^ _zz_151_) ^ _zz_87_[4]) ^ _zz_87_[5]) ^ _zz_87_[6]) ^ _zz_87_[7]) ^ _zz_87_[8]) ^ _zz_87_[9]) ^ _zz_87_[10]) ^ _zz_87_[11]) ^ _zz_87_[12]) ^ _zz_87_[13]) ^ _zz_87_[14]) ^ _zz_87_[15]) ^ _zz_87_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_86_ == io_targetState)))begin
        found[27] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_88_ <= io_startState;
    end
    if(searching)begin
      _zz_88_ <= {_zz_88_[15 : 0],((((((((((((((_zz_152_ ^ _zz_153_) ^ _zz_89_[4]) ^ _zz_89_[5]) ^ _zz_89_[6]) ^ _zz_89_[7]) ^ _zz_89_[8]) ^ _zz_89_[9]) ^ _zz_89_[10]) ^ _zz_89_[11]) ^ _zz_89_[12]) ^ _zz_89_[13]) ^ _zz_89_[14]) ^ _zz_89_[15]) ^ _zz_89_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_88_ == io_targetState)))begin
        found[28] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_90_ <= io_startState;
    end
    if(searching)begin
      _zz_90_ <= {_zz_90_[15 : 0],((((((((((((((_zz_154_ ^ _zz_155_) ^ _zz_91_[4]) ^ _zz_91_[5]) ^ _zz_91_[6]) ^ _zz_91_[7]) ^ _zz_91_[8]) ^ _zz_91_[9]) ^ _zz_91_[10]) ^ _zz_91_[11]) ^ _zz_91_[12]) ^ _zz_91_[13]) ^ _zz_91_[14]) ^ _zz_91_[15]) ^ _zz_91_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_90_ == io_targetState)))begin
        found[29] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_92_ <= io_startState;
    end
    if(searching)begin
      _zz_92_ <= {_zz_92_[15 : 0],((((((((((((((_zz_156_ ^ _zz_157_) ^ _zz_93_[4]) ^ _zz_93_[5]) ^ _zz_93_[6]) ^ _zz_93_[7]) ^ _zz_93_[8]) ^ _zz_93_[9]) ^ _zz_93_[10]) ^ _zz_93_[11]) ^ _zz_93_[12]) ^ _zz_93_[13]) ^ _zz_93_[14]) ^ _zz_93_[15]) ^ _zz_93_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_92_ == io_targetState)))begin
        found[30] <= 1'b1;
        searching <= 1'b0;
      end
    end
    if((io_start_valid && io_start_ready))begin
      _zz_94_ <= io_startState;
    end
    if(searching)begin
      _zz_94_ <= {_zz_94_[15 : 0],((((((((((((((_zz_158_ ^ _zz_159_) ^ _zz_95_[4]) ^ _zz_95_[5]) ^ _zz_95_[6]) ^ _zz_95_[7]) ^ _zz_95_[8]) ^ _zz_95_[9]) ^ _zz_95_[10]) ^ _zz_95_[11]) ^ _zz_95_[12]) ^ _zz_95_[13]) ^ _zz_95_[14]) ^ _zz_95_[15]) ^ _zz_95_[16])};
      if(((counter[9 : 2] == (8'b00000000)) && (_zz_94_ == io_targetState)))begin
        found[31] <= 1'b1;
        searching <= 1'b0;
      end
    end
  end

  always @ (posedge Slow_clk) begin
    searching_regNext <= searching;
  end

endmodule
